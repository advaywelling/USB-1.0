`timescale 1ns / 10ps

module byte_register #(
    // parameters
) (
    input clk, n_rst
);



endmodule

